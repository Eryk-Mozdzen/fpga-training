module project (
    input wire a,
    input wire b,
    output wire y
);

    assign y = a & b; // AND gate

endmodule
